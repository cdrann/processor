`ifndef DEFINE_SV
`define DEFINE_SV
  `define ADDR_BITS 8
  `define DATA_BITS 8
  
  `define OUT 8'h00
  `define SET 8'h01
  `define MOVE 8'h02
  `define JUMP 8'h03
  `define INC 8'h04
  `define DEC 8'h05
  `define SUM 8'h06
  `define SUB 8'h07
  `define MULT 8'h08
  `define DIV 8'h09
  `define AND 8'h0a
  `define OR 8'h0b
  `define XOR 8'h0c
  `define COMP 8'h0d
`endif